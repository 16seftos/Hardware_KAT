module test;
  
  reg clk;
  reg [31:0] pc;
  reg [31:0] inst;
  wire r;
  wire j;
  
  dut dut(
    .clk(clk),
    .pc(pc),
    .inst(inst),
    .r(r),
    .j(j));
  
  initial begin
    //dump waves
    $dumpfile("dump.vcd");
    $dumpvars(1,test);
    clk = 0;
    
   #10 pc = 32'b00001100000000000000000000000000;
       inst = 32'b00001100000000000000000000000001;
   #10 pc = 32'b00011100000000000000000000000000;
       inst = 32'b00000000000000000000000000000000;
   #10 pc = 32'b00111100000000000000000000000000;
       inst = 32'b00000000000110000100000000001000;
   #10 pc = 32'b01011100000000000000000000000000;
       inst = 32'b01000000100000000100000100001100;
   #10 pc = 32'b01011100000000000000000000000000;
       inst = 32'b01000000100110000100000100001100;
    
   #10 $finish;
    
  end
  
  always #5 clk = ~clk;
  
endmodule